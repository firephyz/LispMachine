`ifndef memory_include
`define memory_include

`define memory_data_width 24
`define memory_addr_width 10

`endif