`ifndef alu_include
`define alu_include

`define alu_data_width 16
`define alu_opcode_width 4

`endif