`ifndef memory_include
`define memory_include

`define memory_data_width 24
`define memory_addr_width 10

// Memory unit functions
`define 	GET_CAR			 2'b00
`define 	GET_CDR 			 2'b01
`define 	GET_CONS 		 2'b10
`define 	GET_CONTENTS 	 2'b11

`endif